class Register ;
logic [7:0] data;
static int instance_count = 0;
function new(logic [7:0] value = 8'b0);
    data = value;
    instance_count++;
endfunction

function void load(logic [7:0] value);
    data = value;
endfunction

function logic [7:0] get_data();
    return data;
endfunction

function static int get_instance_count();
    return instance_count;
endfunction

endclass

class shiftLeftRegister extends Register;
    function new(logic [7:0] value = 8'b0);
        super.new(value); 
    endfunction
    
    function void shift_left();
        data = data << 1;
    endfunction
endclass


class shiftRightRegister extends Register;
    function new(logic [7:0] value = 8'b0);
        super.new(value);
    endfunction
    
    function void shift_right();
        this.data = this.data >> 1;
    endfunction
endclass